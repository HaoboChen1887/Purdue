// $Id: $
// File name:   tb_usb_receiver.sv
// Created:     2/22/2018
// Author:      Haobo Chen
// Lab Section: 337-05
// Version:     1.0  Initial Design Entry
// Description: tb_usb_receiver

module tb_usb_receiver();
timeunit 1ns;
	parameter CLK_PERIOD = 64ns;
	reg clk;
	reg clk2;
	reg n_rst;
	reg d_plus;
	reg d_minus;
	reg r_enable;
	reg [7:0]r_data;
	reg empty;
	reg full;
	reg rcving;
	reg r_error;
	usb_receiver TOP(.clk(clk2), .n_rst(n_rst), .d_plus(d_plus), .d_minus(d_minus), .r_enable(r_enable), .r_data(r_data), .empty(empty), .full(full), .rcving(rcving), .r_error(r_error));
	always
	begin
		clk = 1;
		#(CLK_PERIOD / 2);
		clk = 0;
		#(CLK_PERIOD / 2);
	end
	always
	begin
		clk2 = 1;
		#(CLK_PERIOD / 2 / 8);
		clk2 = 0;
		#(CLK_PERIOD / 2 / 8);
	end
	initial
	begin
		//TEST CASE SYNC
		n_rst = 0;
		#(CLK_PERIOD * 5);
		#(CLK_PERIOD * 5);
		r_enable = 0;
		n_rst = 1;	
		d_plus = 1;	
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);	
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);	
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);	
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);	
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);	
		//TEST CASE SHIFT IN + GOOD EOP
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);	
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);	
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);	
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);	
		d_plus = 0;
		d_minus = 0;
		#(CLK_PERIOD);	
		d_plus = 0;
		d_minus = 0;
		#(CLK_PERIOD);	
		d_plus = 1;
		d_minus = 0;
		//TEST 3 SYNC 
		d_plus = 1;	
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);	
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);	
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);	
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);	
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);
		//TEST 4
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);	
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 0;
		d_minus = 0;
		#(CLK_PERIOD);	
		d_plus = 0;
		d_minus = 0;
		#(CLK_PERIOD);	
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);
		//TEST 5 SYNC
		d_plus = 1;	
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);	
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);	
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);	
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);	
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);
		//PACKET1
		d_plus = 1;	
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);	
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);	
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);	
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);	
		r_enable = 1;
		#(CLK_PERIOD);
		r_enable = 0;
		//PACKET2
		d_plus = 1;	
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);	
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);	
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);	
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);
		r_enable = 1;
		#(CLK_PERIOD);
		r_enable = 0;
		//PACKET3
		d_plus = 1;	
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);	
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);	
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);	
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);	
		//EOP
		d_plus = 0;
		d_minus = 0;
		#(CLK_PERIOD);	
		d_plus = 0;
		d_minus = 0;
		#(CLK_PERIOD);	
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);
		//TEST 6
		d_plus = 1;	
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);	
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);	
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);	
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);	
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);
		//PACKET1
		d_plus = 0;	
		d_minus = 1;
		#(CLK_PERIOD);
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);	
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);	
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);	
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);	
		//PACKET2
		d_plus = 0;	
		d_minus = 1;
		#(CLK_PERIOD);
		d_plus = 0;
		d_minus = 1;
		#(CLK_PERIOD);
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);
		//EOP	
		d_plus = 0;
		d_minus = 0;
		#(CLK_PERIOD);	
		d_plus = 0;
		d_minus = 0;
		#(CLK_PERIOD);	
		d_plus = 1;
		d_minus = 0;
		#(CLK_PERIOD);
	end
endmodule

